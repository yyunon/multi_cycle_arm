module PC #(parameter W=32)(input )